// Global nets module 

`celldefine
module cds_globals;


wire VDD_;


endmodule
`endcelldefine
